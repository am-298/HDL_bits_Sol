////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////
// 
// implementation of ground  module
//
////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////


module top_module (
    output out);
    
    assign out = 1'b0;

endmodule
