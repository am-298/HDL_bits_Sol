
////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////
// Author : Ayushi Maurya
//// wire type connection example
//
////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////
module top_module (
    input in,
    output out);
    
    wire out1=in;
    
    assign out = out1 ;

endmodule